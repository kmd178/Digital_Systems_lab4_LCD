`timescale 1ns / 1ps
module lcd_controller(




    );


endmodule
